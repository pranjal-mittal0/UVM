/*-----------------------------------------------------------------
File name     : packet_pkg.sv
Developers    : Pranjal Mittal
Created       : 25/05/2023
Description   : lab3 packet data item 
Notes         : From the Cadence "Essential SystemVerilog for UVM" training
-------------------------------------------------------------------
This is for lab work for the above training.

-----------------------------------------------------------------*/
package packet_pkg;
    `include "packet_data.sv"
endpackage