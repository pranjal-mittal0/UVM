/*-----------------------------------------------------------------
File name     : sequence_item.sv
Developers    : Pranjal Mittal
Created       : 12/05/2023
Description   : 
-------------------------------------------------------------------*/