/*-----------------------------------------------------------------
File name     : sequencer.sv
Developers    : Pranjal Mittal
Created       : 30/05/2023
Description   : lab6 sequencer class
Notes         : From the Cadence "Essential SystemVerilog for UVM" training
-------------------------------------------------------------------
This is for lab work for the above training.

-----------------------------------------------------------------*/
class sequencer extends component_base;
    int portno; //will be set in configuration and used to assign source for packets generated by sequencer.
    int ok;
    function new(string name,component_base parent);
        super.new(name,parent);
    endfunction //new()

    function void get_next_item(output packet pkt);
        //packet pkt; //already declared in the argument.
        psingle ps;
        pmulticast pm;
        pbroadcast pb;
        randcase
            1:begin : single_packet
                ps=new("ps",portno);
                ok=ps.randomize();
                pkt=ps;
            end
            1:begin : multicast_packet
                pm=new("pm",portno);
                ok=pm.randomize();
                pkt=pm;
            end
            1: begin : broadcast_packet
                pb=new("pb",portno);
                ok=pb.randomize();
                pkt=pb;
            end
        endcase
    endfunction
endclass //sequencer extends component_base