/*-----------------------------------------------------------------
File name     : sequence.sv
Developers    : Pranjal Mittal
Created       : 12/05/2023
Description   : 
-------------------------------------------------------------------*/