/*-----------------------------------------------------------------
File name     : packet_p.sv
Developers    : Brian Dickinson
Created       : 01/08/19
Description   : lab4 packet data package
Notes         : From the Cadence "Essential SystemVerilog for UVM" training
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2019
-----------------------------------------------------------------*/

package packet_pkg;

`include "packet_data.sv"

endpackage
